`timescale 1ns / 1ps
module PCAdder(
	input  Pc,
	output PCPlus
    );
	 assign pCPlus = Pc + 4;


endmodule
