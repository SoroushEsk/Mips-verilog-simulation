`timescale 1ns / 1ps

module IFIDRegister(
    );


endmodule
